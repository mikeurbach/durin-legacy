module f(x);
   output[63:0] x;

   assign x = 2+2;
   
endmodule // f
